magic
tech scmos
timestamp 1666954522
<< pwell >>
rect -8 -10 11 5
<< nwell >>
rect -8 12 11 27
<< polysilicon >>
rect 0 16 2 18
rect 0 10 2 13
rect 0 3 2 6
rect 0 -2 2 0
<< ndiffusion >>
rect -1 0 0 3
rect 2 0 4 3
<< pdiffusion >>
rect -1 13 0 16
rect 2 13 4 16
<< metal1 >>
rect -1 21 3 25
rect -5 17 -2 21
rect 5 10 8 13
rect -6 6 -2 10
rect 5 7 9 10
rect 5 3 8 7
rect -5 -5 -2 -1
rect -1 -9 3 -5
<< ntransistor >>
rect 0 0 2 3
<< ptransistor >>
rect 0 13 2 16
<< polycontact >>
rect -2 6 2 10
<< ndcontact >>
rect -5 -1 -1 3
rect 4 -1 8 3
<< pdcontact >>
rect -5 13 -1 17
rect 4 13 8 17
<< psubstratepcontact >>
rect -5 -9 -1 -5
rect 3 -9 7 -5
<< nsubstratencontact >>
rect -5 21 -1 25
rect 3 21 7 25
<< labels >>
rlabel metal1 1 23 1 23 5 vdd!
rlabel metal1 1 -7 1 -7 1 gnd!
rlabel metal1 -6 6 -6 10 3 in
rlabel metal1 9 7 9 10 7 out
<< end >>
