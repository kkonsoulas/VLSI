*
.include MOSIS_TSMC_025um.spice


.option scale=1u


MNMOS1 out1 in vdd 0 CMOSN w=3 l=2


Cout2 out1 0 0.1pF

vvdd vdd 0 2.5V DC
vgs in 0 2.5V  DC
* vvdd vdd 0 2.5 DC
.ic V(out1)=0V
* .ic V(out1)=0

.tran 100ns 1ms
* .plot dc v(out)

.control
    run
    meas tran volout1 
    + find v(out1) at=1ms
    plot v(out1) title "Voltage drop for one NMOS"
.endc



.end

