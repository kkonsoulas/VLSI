magic
tech scmos
timestamp 1670351680
<< pwell >>
rect -11 -22 25 -2
<< nwell >>
rect -11 17 25 48
<< polysilicon >>
rect -6 48 -4 50
rect 2 48 4 50
rect 10 48 12 50
rect 18 28 20 30
rect -6 -6 -4 18
rect 2 8 4 18
rect 10 8 12 18
rect 18 8 20 18
rect 3 4 4 8
rect 11 4 12 8
rect 19 4 20 8
rect 2 -6 4 4
rect 10 -6 12 4
rect 18 -6 20 4
rect -6 -16 -4 -14
rect 2 -16 4 -14
rect 10 -16 12 -14
rect 18 -16 20 -14
<< ndiffusion >>
rect -7 -14 -6 -6
rect -4 -14 -3 -6
rect 1 -14 2 -6
rect 4 -14 5 -6
rect 9 -14 10 -6
rect 12 -14 13 -6
rect 17 -14 18 -6
rect 20 -14 21 -6
<< pdiffusion >>
rect -7 18 -6 48
rect -4 18 2 48
rect 4 18 10 48
rect 12 18 13 48
rect 17 18 18 28
rect 20 18 21 28
<< metal1 >>
rect -11 51 25 54
rect -11 48 -7 51
rect 21 48 25 51
rect 21 28 25 32
rect 13 15 17 18
rect 13 12 25 15
rect -11 4 -10 8
rect -2 4 -1 8
rect 6 4 7 8
rect 14 4 15 8
rect -3 -3 17 0
rect -3 -6 1 -3
rect 13 -6 17 -3
rect 22 -6 25 12
rect -11 -18 -7 -14
rect 5 -18 9 -14
<< ntransistor >>
rect -6 -14 -4 -6
rect 2 -14 4 -6
rect 10 -14 12 -6
rect 18 -14 20 -6
<< ptransistor >>
rect -6 18 -4 48
rect 2 18 4 48
rect 10 18 12 48
rect 18 18 20 28
<< polycontact >>
rect -10 4 -6 8
rect -1 4 3 8
rect 7 4 11 8
rect 15 4 19 8
<< ndcontact >>
rect -11 -14 -7 -6
rect -3 -14 1 -6
rect 5 -14 9 -6
rect 13 -14 17 -6
rect 21 -14 25 -6
<< pdcontact >>
rect -11 18 -7 48
rect 13 18 17 48
rect 21 18 25 28
<< psubstratepcontact >>
rect -11 -22 25 -18
<< nsubstratencontact >>
rect 21 32 25 48
<< labels >>
rlabel psubstratepcontact -11 -22 -11 -18 2 gnd
rlabel metal1 25 -6 25 15 7 out
rlabel metal1 -11 4 -11 8 3 a
rlabel metal1 -2 4 -2 8 1 c
rlabel metal1 6 4 6 8 1 d
rlabel metal1 14 4 14 8 1 b
rlabel nsubstratencontact 25 32 25 48 7 Vdd
<< end >>
